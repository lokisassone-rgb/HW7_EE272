../results/conv.lef